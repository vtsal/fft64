library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity realcoeff64 is
    generic(SIZE: integer;
	        WIDTH: integer:=18);
	port(
        index 		: in  std_logic_vector(2*SIZE-2 downto 0);
        coeff 		: out std_logic_vector(WIDTH-1 downto 0)
    );
end realcoeff64;

ARCHITECTURE dataflow OF realcoeff64 IS

SIGNAL indx: INTEGER RANGE 0 TO (2**SIZE)*(2**(SIZE-1))-1;
TYPE vector_array IS ARRAY (0 to (2**SIZE)*(2**(SIZE-1))-1) OF STD_LOGIC_VECTOR(((WIDTH+4-1)/4)*4-1 DOWNTO 0);
CONSTANT memory : vector_array := 
	(

--64 point FFT coefficients
--Row 0
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
--Row 1
x"00400",
x"3fc00",
x"00000",
x"00000",
x"002d4",
x"3fd2c",
x"3fd2c",
x"002d4",
x"003b2",
x"3fc4e",
x"3fcf1",
x"0030f",
x"0030f",
x"3fcf1",
x"3fc4e",
x"003b2",
x"003ec",
x"3fc14",
x"3fce1",
x"0031f",
x"00238",
x"3fdc8",
x"3fcad",
x"00353",
x"00353",
x"3fcad",
x"3fdc8",
x"00238",
x"0031f",
x"3fce1",
x"3fc14",
x"003ec",
x"003fb",
x"3fc05",
x"3fcde",
x"00322",
x"00289",
x"3fd77",
x"3fce9",
x"00317",
x"00387",
x"3fc79",
x"3fc3b",
x"003c5",
x"00252",
x"3fdae",
x"3fc2d",
x"003d3",
x"003d3",
x"3fc2d",
x"3fdae",
x"00252",
x"003c5",
x"3fc3b",
x"3fc79",
x"00387",
x"00317",
x"3fce9",
x"3fd77",
x"00289",
x"00322",
x"3fcde",
x"3fc05",
x"003fb",
--Row 2
x"00400",
x"00400",
x"3fc00",
x"3fc00",
x"00000",
x"00000",
x"00000",
x"00000",
x"002d4",
x"002d4",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"002d4",
x"002d4",
x"003b2",
x"003b2",
x"3fc4e",
x"3fc4e",
x"3fcf1",
x"3fcf1",
x"0030f",
x"0030f",
x"0030f",
x"0030f",
x"3fcf1",
x"3fcf1",
x"3fc4e",
x"3fc4e",
x"003b2",
x"003b2",
x"003ec",
x"003ec",
x"3fc14",
x"3fc14",
x"3fce1",
x"3fce1",
x"0031f",
x"0031f",
x"00238",
x"00238",
x"3fdc8",
x"3fdc8",
x"3fcad",
x"3fcad",
x"00353",
x"00353",
x"00353",
x"00353",
x"3fcad",
x"3fcad",
x"3fdc8",
x"3fdc8",
x"00238",
x"00238",
x"0031f",
x"0031f",
x"3fce1",
x"3fce1",
x"3fc14",
x"3fc14",
x"003ec",
x"003ec",
--Row 3
x"00400",
x"3fc00",
x"00000",
x"00000",
x"3fd2c",
x"002d4",
x"002d4",
x"3fd2c",
x"0030f",
x"3fcf1",
x"003b2",
x"3fc4e",
x"3fc4e",
x"003b2",
x"3fcf1",
x"0030f",
x"00353",
x"3fcad",
x"00238",
x"3fdc8",
x"3fc14",
x"003ec",
x"0031f",
x"3fce1",
x"3fce1",
x"0031f",
x"003ec",
x"3fc14",
x"3fdc8",
x"00238",
x"3fcad",
x"00353",
x"003d3",
x"3fc2d",
x"00252",
x"3fdae",
x"3fc79",
x"00387",
x"003c5",
x"3fc3b",
x"00322",
x"3fcde",
x"003fb",
x"3fc05",
x"3fce9",
x"00317",
x"3fd77",
x"00289",
x"00289",
x"3fd77",
x"00317",
x"3fce9",
x"3fc05",
x"003fb",
x"3fcde",
x"00322",
x"3fc3b",
x"003c5",
x"00387",
x"3fc79",
x"3fdae",
x"00252",
x"3fc2d",
x"003d3",
--Row 4
x"00400",
x"00400",
x"00400",
x"00400",
x"3fc00",
x"3fc00",
x"3fc00",
x"3fc00",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"002d4",
x"002d4",
x"002d4",
x"002d4",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"002d4",
x"002d4",
x"002d4",
x"002d4",
x"003b2",
x"003b2",
x"003b2",
x"003b2",
x"3fc4e",
x"3fc4e",
x"3fc4e",
x"3fc4e",
x"3fcf1",
x"3fcf1",
x"3fcf1",
x"3fcf1",
x"0030f",
x"0030f",
x"0030f",
x"0030f",
x"0030f",
x"0030f",
x"0030f",
x"0030f",
x"3fcf1",
x"3fcf1",
x"3fcf1",
x"3fcf1",
x"3fc4e",
x"3fc4e",
x"3fc4e",
x"3fc4e",
x"003b2",
x"003b2",
x"003b2",
x"003b2",
--Row 5
x"00400",
x"3fc00",
x"00000",
x"00000",
x"3fd2c",
x"002d4",
x"002d4",
x"3fd2c",
x"3fcf1",
x"0030f",
x"3fc4e",
x"003b2",
x"003b2",
x"3fc4e",
x"0030f",
x"3fcf1",
x"00238",
x"3fdc8",
x"3fcad",
x"00353",
x"0031f",
x"3fce1",
x"003ec",
x"3fc14",
x"3fc14",
x"003ec",
x"3fce1",
x"0031f",
x"00353",
x"3fcad",
x"3fdc8",
x"00238",
x"00387",
x"3fc79",
x"3fc3b",
x"003c5",
x"3fdae",
x"00252",
x"003d3",
x"3fc2d",
x"3fce9",
x"00317",
x"3fd77",
x"00289",
x"003fb",
x"3fc05",
x"3fcde",
x"00322",
x"00322",
x"3fcde",
x"3fc05",
x"003fb",
x"00289",
x"3fd77",
x"00317",
x"3fce9",
x"3fc2d",
x"003d3",
x"00252",
x"3fdae",
x"003c5",
x"3fc3b",
x"3fc79",
x"00387",
--Row 6
x"00400",
x"00400",
x"3fc00",
x"3fc00",
x"00000",
x"00000",
x"00000",
x"00000",
x"3fd2c",
x"3fd2c",
x"002d4",
x"002d4",
x"002d4",
x"002d4",
x"3fd2c",
x"3fd2c",
x"0030f",
x"0030f",
x"3fcf1",
x"3fcf1",
x"003b2",
x"003b2",
x"3fc4e",
x"3fc4e",
x"3fc4e",
x"3fc4e",
x"003b2",
x"003b2",
x"3fcf1",
x"3fcf1",
x"0030f",
x"0030f",
x"00353",
x"00353",
x"3fcad",
x"3fcad",
x"00238",
x"00238",
x"3fdc8",
x"3fdc8",
x"3fc14",
x"3fc14",
x"003ec",
x"003ec",
x"0031f",
x"0031f",
x"3fce1",
x"3fce1",
x"3fce1",
x"3fce1",
x"0031f",
x"0031f",
x"003ec",
x"003ec",
x"3fc14",
x"3fc14",
x"3fdc8",
x"3fdc8",
x"00238",
x"00238",
x"3fcad",
x"3fcad",
x"00353",
x"00353",
--Row 7
x"00400",
x"3fc00",
x"00000",
x"00000",
x"002d4",
x"3fd2c",
x"3fd2c",
x"002d4",
x"3fc4e",
x"003b2",
x"0030f",
x"3fcf1",
x"3fcf1",
x"0030f",
x"003b2",
x"3fc4e",
x"0031f",
x"3fce1",
x"003ec",
x"3fc14",
x"00353",
x"3fcad",
x"00238",
x"3fdc8",
x"3fdc8",
x"00238",
x"3fcad",
x"00353",
x"3fc14",
x"003ec",
x"3fce1",
x"0031f",
x"00317",
x"3fce9",
x"00289",
x"3fd77",
x"003fb",
x"3fc05",
x"3fcde",
x"00322",
x"3fc2d",
x"003d3",
x"3fdae",
x"00252",
x"3fc79",
x"00387",
x"003c5",
x"3fc3b",
x"3fc3b",
x"003c5",
x"00387",
x"3fc79",
x"00252",
x"3fdae",
x"003d3",
x"3fc2d",
x"00322",
x"3fcde",
x"3fc05",
x"003fb",
x"3fd77",
x"00289",
x"3fce9",
x"00317",
--Row 8
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"3fc00",
x"3fc00",
x"3fc00",
x"3fc00",
x"3fc00",
x"3fc00",
x"3fc00",
x"3fc00",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"002d4",
x"002d4",
x"002d4",
x"002d4",
x"002d4",
x"002d4",
x"002d4",
x"002d4",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"002d4",
x"002d4",
x"002d4",
x"002d4",
x"002d4",
x"002d4",
x"002d4",
x"002d4",
--Row 9
x"00400",
x"3fc00",
x"00000",
x"00000",
x"002d4",
x"3fd2c",
x"3fd2c",
x"002d4",
x"3fc4e",
x"003b2",
x"0030f",
x"3fcf1",
x"3fcf1",
x"0030f",
x"003b2",
x"3fc4e",
x"3fce1",
x"0031f",
x"3fc14",
x"003ec",
x"3fcad",
x"00353",
x"3fdc8",
x"00238",
x"00238",
x"3fdc8",
x"00353",
x"3fcad",
x"003ec",
x"3fc14",
x"0031f",
x"3fce1",
x"00289",
x"3fd77",
x"3fce9",
x"00317",
x"3fcde",
x"00322",
x"3fc05",
x"003fb",
x"3fdae",
x"00252",
x"003d3",
x"3fc2d",
x"003c5",
x"3fc3b",
x"00387",
x"3fc79",
x"3fc79",
x"00387",
x"3fc3b",
x"003c5",
x"3fc2d",
x"003d3",
x"00252",
x"3fdae",
x"003fb",
x"3fc05",
x"00322",
x"3fcde",
x"00317",
x"3fce9",
x"3fd77",
x"00289",
--Row 10
x"00400",
x"00400",
x"3fc00",
x"3fc00",
x"00000",
x"00000",
x"00000",
x"00000",
x"3fd2c",
x"3fd2c",
x"002d4",
x"002d4",
x"002d4",
x"002d4",
x"3fd2c",
x"3fd2c",
x"3fcf1",
x"3fcf1",
x"0030f",
x"0030f",
x"3fc4e",
x"3fc4e",
x"003b2",
x"003b2",
x"003b2",
x"003b2",
x"3fc4e",
x"3fc4e",
x"0030f",
x"0030f",
x"3fcf1",
x"3fcf1",
x"00238",
x"00238",
x"3fdc8",
x"3fdc8",
x"3fcad",
x"3fcad",
x"00353",
x"00353",
x"0031f",
x"0031f",
x"3fce1",
x"3fce1",
x"003ec",
x"003ec",
x"3fc14",
x"3fc14",
x"3fc14",
x"3fc14",
x"003ec",
x"003ec",
x"3fce1",
x"3fce1",
x"0031f",
x"0031f",
x"00353",
x"00353",
x"3fcad",
x"3fcad",
x"3fdc8",
x"3fdc8",
x"00238",
x"00238",
--Row 11
x"00400",
x"3fc00",
x"00000",
x"00000",
x"3fd2c",
x"002d4",
x"002d4",
x"3fd2c",
x"3fcf1",
x"0030f",
x"3fc4e",
x"003b2",
x"003b2",
x"3fc4e",
x"0030f",
x"3fcf1",
x"3fdc8",
x"00238",
x"00353",
x"3fcad",
x"3fce1",
x"0031f",
x"3fc14",
x"003ec",
x"003ec",
x"3fc14",
x"0031f",
x"3fce1",
x"3fcad",
x"00353",
x"00238",
x"3fdc8",
x"003c5",
x"3fc3b",
x"00387",
x"3fc79",
x"3fc2d",
x"003d3",
x"3fdae",
x"00252",
x"00289",
x"3fd77",
x"3fce9",
x"00317",
x"00322",
x"3fcde",
x"003fb",
x"3fc05",
x"3fc05",
x"003fb",
x"3fcde",
x"00322",
x"00317",
x"3fce9",
x"3fd77",
x"00289",
x"00252",
x"3fdae",
x"003d3",
x"3fc2d",
x"3fc79",
x"00387",
x"3fc3b",
x"003c5",
--Row 12
x"00400",
x"00400",
x"00400",
x"00400",
x"3fc00",
x"3fc00",
x"3fc00",
x"3fc00",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"002d4",
x"002d4",
x"002d4",
x"002d4",
x"002d4",
x"002d4",
x"002d4",
x"002d4",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"0030f",
x"0030f",
x"0030f",
x"0030f",
x"3fcf1",
x"3fcf1",
x"3fcf1",
x"3fcf1",
x"003b2",
x"003b2",
x"003b2",
x"003b2",
x"3fc4e",
x"3fc4e",
x"3fc4e",
x"3fc4e",
x"3fc4e",
x"3fc4e",
x"3fc4e",
x"3fc4e",
x"003b2",
x"003b2",
x"003b2",
x"003b2",
x"3fcf1",
x"3fcf1",
x"3fcf1",
x"3fcf1",
x"0030f",
x"0030f",
x"0030f",
x"0030f",
--Row 13
x"00400",
x"3fc00",
x"00000",
x"00000",
x"3fd2c",
x"002d4",
x"002d4",
x"3fd2c",
x"0030f",
x"3fcf1",
x"003b2",
x"3fc4e",
x"3fc4e",
x"003b2",
x"3fcf1",
x"0030f",
x"3fcad",
x"00353",
x"3fdc8",
x"00238",
x"003ec",
x"3fc14",
x"3fce1",
x"0031f",
x"0031f",
x"3fce1",
x"3fc14",
x"003ec",
x"00238",
x"3fdc8",
x"00353",
x"3fcad",
x"00252",
x"3fdae",
x"3fc2d",
x"003d3",
x"003c5",
x"3fc3b",
x"00387",
x"3fc79",
x"003fb",
x"3fc05",
x"3fcde",
x"00322",
x"3fd77",
x"00289",
x"00317",
x"3fce9",
x"3fce9",
x"00317",
x"00289",
x"3fd77",
x"00322",
x"3fcde",
x"3fc05",
x"003fb",
x"3fc79",
x"00387",
x"3fc3b",
x"003c5",
x"003d3",
x"3fc2d",
x"3fdae",
x"00252",
--Row 14
x"00400",
x"00400",
x"3fc00",
x"3fc00",
x"00000",
x"00000",
x"00000",
x"00000",
x"002d4",
x"002d4",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"002d4",
x"002d4",
x"3fc4e",
x"3fc4e",
x"003b2",
x"003b2",
x"0030f",
x"0030f",
x"3fcf1",
x"3fcf1",
x"3fcf1",
x"3fcf1",
x"0030f",
x"0030f",
x"003b2",
x"003b2",
x"3fc4e",
x"3fc4e",
x"0031f",
x"0031f",
x"3fce1",
x"3fce1",
x"003ec",
x"003ec",
x"3fc14",
x"3fc14",
x"00353",
x"00353",
x"3fcad",
x"3fcad",
x"00238",
x"00238",
x"3fdc8",
x"3fdc8",
x"3fdc8",
x"3fdc8",
x"00238",
x"00238",
x"3fcad",
x"3fcad",
x"00353",
x"00353",
x"3fc14",
x"3fc14",
x"003ec",
x"003ec",
x"3fce1",
x"3fce1",
x"0031f",
x"0031f",
--Row 15
x"00400",
x"3fc00",
x"00000",
x"00000",
x"002d4",
x"3fd2c",
x"3fd2c",
x"002d4",
x"003b2",
x"3fc4e",
x"3fcf1",
x"0030f",
x"0030f",
x"3fcf1",
x"3fc4e",
x"003b2",
x"3fc14",
x"003ec",
x"0031f",
x"3fce1",
x"3fdc8",
x"00238",
x"00353",
x"3fcad",
x"3fcad",
x"00353",
x"00238",
x"3fdc8",
x"3fce1",
x"0031f",
x"003ec",
x"3fc14",
x"00322",
x"3fcde",
x"003fb",
x"3fc05",
x"00317",
x"3fce9",
x"00289",
x"3fd77",
x"003c5",
x"3fc3b",
x"00387",
x"3fc79",
x"003d3",
x"3fc2d",
x"00252",
x"3fdae",
x"3fdae",
x"00252",
x"3fc2d",
x"003d3",
x"3fc79",
x"00387",
x"3fc3b",
x"003c5",
x"3fd77",
x"00289",
x"3fce9",
x"00317",
x"3fc05",
x"003fb",
x"3fcde",
x"00322",
--Row 16
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"3fc00",
x"3fc00",
x"3fc00",
x"3fc00",
x"3fc00",
x"3fc00",
x"3fc00",
x"3fc00",
x"3fc00",
x"3fc00",
x"3fc00",
x"3fc00",
x"3fc00",
x"3fc00",
x"3fc00",
x"3fc00",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
--Row 17
x"00400",
x"3fc00",
x"00000",
x"00000",
x"002d4",
x"3fd2c",
x"3fd2c",
x"002d4",
x"003b2",
x"3fc4e",
x"3fcf1",
x"0030f",
x"0030f",
x"3fcf1",
x"3fc4e",
x"003b2",
x"3fc14",
x"003ec",
x"0031f",
x"3fce1",
x"3fdc8",
x"00238",
x"00353",
x"3fcad",
x"3fcad",
x"00353",
x"00238",
x"3fdc8",
x"3fce1",
x"0031f",
x"003ec",
x"3fc14",
x"3fcde",
x"00322",
x"3fc05",
x"003fb",
x"3fce9",
x"00317",
x"3fd77",
x"00289",
x"3fc3b",
x"003c5",
x"3fc79",
x"00387",
x"3fc2d",
x"003d3",
x"3fdae",
x"00252",
x"00252",
x"3fdae",
x"003d3",
x"3fc2d",
x"00387",
x"3fc79",
x"003c5",
x"3fc3b",
x"00289",
x"3fd77",
x"00317",
x"3fce9",
x"003fb",
x"3fc05",
x"00322",
x"3fcde",
--Row 18
x"00400",
x"00400",
x"3fc00",
x"3fc00",
x"00000",
x"00000",
x"00000",
x"00000",
x"002d4",
x"002d4",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"002d4",
x"002d4",
x"3fc4e",
x"3fc4e",
x"003b2",
x"003b2",
x"0030f",
x"0030f",
x"3fcf1",
x"3fcf1",
x"3fcf1",
x"3fcf1",
x"0030f",
x"0030f",
x"003b2",
x"003b2",
x"3fc4e",
x"3fc4e",
x"3fce1",
x"3fce1",
x"0031f",
x"0031f",
x"3fc14",
x"3fc14",
x"003ec",
x"003ec",
x"3fcad",
x"3fcad",
x"00353",
x"00353",
x"3fdc8",
x"3fdc8",
x"00238",
x"00238",
x"00238",
x"00238",
x"3fdc8",
x"3fdc8",
x"00353",
x"00353",
x"3fcad",
x"3fcad",
x"003ec",
x"003ec",
x"3fc14",
x"3fc14",
x"0031f",
x"0031f",
x"3fce1",
x"3fce1",
--Row 19
x"00400",
x"3fc00",
x"00000",
x"00000",
x"3fd2c",
x"002d4",
x"002d4",
x"3fd2c",
x"0030f",
x"3fcf1",
x"003b2",
x"3fc4e",
x"3fc4e",
x"003b2",
x"3fcf1",
x"0030f",
x"3fcad",
x"00353",
x"3fdc8",
x"00238",
x"003ec",
x"3fc14",
x"3fce1",
x"0031f",
x"0031f",
x"3fce1",
x"3fc14",
x"003ec",
x"00238",
x"3fdc8",
x"00353",
x"3fcad",
x"3fdae",
x"00252",
x"003d3",
x"3fc2d",
x"3fc3b",
x"003c5",
x"3fc79",
x"00387",
x"3fc05",
x"003fb",
x"00322",
x"3fcde",
x"00289",
x"3fd77",
x"3fce9",
x"00317",
x"00317",
x"3fce9",
x"3fd77",
x"00289",
x"3fcde",
x"00322",
x"003fb",
x"3fc05",
x"00387",
x"3fc79",
x"003c5",
x"3fc3b",
x"3fc2d",
x"003d3",
x"00252",
x"3fdae",
--Row 20
x"00400",
x"00400",
x"00400",
x"00400",
x"3fc00",
x"3fc00",
x"3fc00",
x"3fc00",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"002d4",
x"002d4",
x"002d4",
x"002d4",
x"002d4",
x"002d4",
x"002d4",
x"002d4",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"3fcf1",
x"3fcf1",
x"3fcf1",
x"3fcf1",
x"0030f",
x"0030f",
x"0030f",
x"0030f",
x"3fc4e",
x"3fc4e",
x"3fc4e",
x"3fc4e",
x"003b2",
x"003b2",
x"003b2",
x"003b2",
x"003b2",
x"003b2",
x"003b2",
x"003b2",
x"3fc4e",
x"3fc4e",
x"3fc4e",
x"3fc4e",
x"0030f",
x"0030f",
x"0030f",
x"0030f",
x"3fcf1",
x"3fcf1",
x"3fcf1",
x"3fcf1",
--Row 21
x"00400",
x"3fc00",
x"00000",
x"00000",
x"3fd2c",
x"002d4",
x"002d4",
x"3fd2c",
x"3fcf1",
x"0030f",
x"3fc4e",
x"003b2",
x"003b2",
x"3fc4e",
x"0030f",
x"3fcf1",
x"3fdc8",
x"00238",
x"00353",
x"3fcad",
x"3fce1",
x"0031f",
x"3fc14",
x"003ec",
x"003ec",
x"3fc14",
x"0031f",
x"3fce1",
x"3fcad",
x"00353",
x"00238",
x"3fdc8",
x"3fc3b",
x"003c5",
x"3fc79",
x"00387",
x"003d3",
x"3fc2d",
x"00252",
x"3fdae",
x"3fd77",
x"00289",
x"00317",
x"3fce9",
x"3fcde",
x"00322",
x"3fc05",
x"003fb",
x"003fb",
x"3fc05",
x"00322",
x"3fcde",
x"3fce9",
x"00317",
x"00289",
x"3fd77",
x"3fdae",
x"00252",
x"3fc2d",
x"003d3",
x"00387",
x"3fc79",
x"003c5",
x"3fc3b",
--Row 22
x"00400",
x"00400",
x"3fc00",
x"3fc00",
x"00000",
x"00000",
x"00000",
x"00000",
x"3fd2c",
x"3fd2c",
x"002d4",
x"002d4",
x"002d4",
x"002d4",
x"3fd2c",
x"3fd2c",
x"3fcf1",
x"3fcf1",
x"0030f",
x"0030f",
x"3fc4e",
x"3fc4e",
x"003b2",
x"003b2",
x"003b2",
x"003b2",
x"3fc4e",
x"3fc4e",
x"0030f",
x"0030f",
x"3fcf1",
x"3fcf1",
x"3fdc8",
x"3fdc8",
x"00238",
x"00238",
x"00353",
x"00353",
x"3fcad",
x"3fcad",
x"3fce1",
x"3fce1",
x"0031f",
x"0031f",
x"3fc14",
x"3fc14",
x"003ec",
x"003ec",
x"003ec",
x"003ec",
x"3fc14",
x"3fc14",
x"0031f",
x"0031f",
x"3fce1",
x"3fce1",
x"3fcad",
x"3fcad",
x"00353",
x"00353",
x"00238",
x"00238",
x"3fdc8",
x"3fdc8",
--Row 23
x"00400",
x"3fc00",
x"00000",
x"00000",
x"002d4",
x"3fd2c",
x"3fd2c",
x"002d4",
x"3fc4e",
x"003b2",
x"0030f",
x"3fcf1",
x"3fcf1",
x"0030f",
x"003b2",
x"3fc4e",
x"3fce1",
x"0031f",
x"3fc14",
x"003ec",
x"3fcad",
x"00353",
x"3fdc8",
x"00238",
x"00238",
x"3fdc8",
x"00353",
x"3fcad",
x"003ec",
x"3fc14",
x"0031f",
x"3fce1",
x"3fd77",
x"00289",
x"00317",
x"3fce9",
x"00322",
x"3fcde",
x"003fb",
x"3fc05",
x"00252",
x"3fdae",
x"3fc2d",
x"003d3",
x"3fc3b",
x"003c5",
x"3fc79",
x"00387",
x"00387",
x"3fc79",
x"003c5",
x"3fc3b",
x"003d3",
x"3fc2d",
x"3fdae",
x"00252",
x"3fc05",
x"003fb",
x"3fcde",
x"00322",
x"3fce9",
x"00317",
x"00289",
x"3fd77",
--Row 24
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"00400",
x"3fc00",
x"3fc00",
x"3fc00",
x"3fc00",
x"3fc00",
x"3fc00",
x"3fc00",
x"3fc00",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"002d4",
x"002d4",
x"002d4",
x"002d4",
x"002d4",
x"002d4",
x"002d4",
x"002d4",
x"002d4",
x"002d4",
x"002d4",
x"002d4",
x"002d4",
x"002d4",
x"002d4",
x"002d4",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"3fd2c",
--Row 25
x"00400",
x"3fc00",
x"00000",
x"00000",
x"002d4",
x"3fd2c",
x"3fd2c",
x"002d4",
x"3fc4e",
x"003b2",
x"0030f",
x"3fcf1",
x"3fcf1",
x"0030f",
x"003b2",
x"3fc4e",
x"0031f",
x"3fce1",
x"003ec",
x"3fc14",
x"00353",
x"3fcad",
x"00238",
x"3fdc8",
x"3fdc8",
x"00238",
x"3fcad",
x"00353",
x"3fc14",
x"003ec",
x"3fce1",
x"0031f",
x"3fce9",
x"00317",
x"3fd77",
x"00289",
x"3fc05",
x"003fb",
x"00322",
x"3fcde",
x"003d3",
x"3fc2d",
x"00252",
x"3fdae",
x"00387",
x"3fc79",
x"3fc3b",
x"003c5",
x"003c5",
x"3fc3b",
x"3fc79",
x"00387",
x"3fdae",
x"00252",
x"3fc2d",
x"003d3",
x"3fcde",
x"00322",
x"003fb",
x"3fc05",
x"00289",
x"3fd77",
x"00317",
x"3fce9",
--Row 26
x"00400",
x"00400",
x"3fc00",
x"3fc00",
x"00000",
x"00000",
x"00000",
x"00000",
x"3fd2c",
x"3fd2c",
x"002d4",
x"002d4",
x"002d4",
x"002d4",
x"3fd2c",
x"3fd2c",
x"0030f",
x"0030f",
x"3fcf1",
x"3fcf1",
x"003b2",
x"003b2",
x"3fc4e",
x"3fc4e",
x"3fc4e",
x"3fc4e",
x"003b2",
x"003b2",
x"3fcf1",
x"3fcf1",
x"0030f",
x"0030f",
x"3fcad",
x"3fcad",
x"00353",
x"00353",
x"3fdc8",
x"3fdc8",
x"00238",
x"00238",
x"003ec",
x"003ec",
x"3fc14",
x"3fc14",
x"3fce1",
x"3fce1",
x"0031f",
x"0031f",
x"0031f",
x"0031f",
x"3fce1",
x"3fce1",
x"3fc14",
x"3fc14",
x"003ec",
x"003ec",
x"00238",
x"00238",
x"3fdc8",
x"3fdc8",
x"00353",
x"00353",
x"3fcad",
x"3fcad",
--Row 27
x"00400",
x"3fc00",
x"00000",
x"00000",
x"3fd2c",
x"002d4",
x"002d4",
x"3fd2c",
x"3fcf1",
x"0030f",
x"3fc4e",
x"003b2",
x"003b2",
x"3fc4e",
x"0030f",
x"3fcf1",
x"00238",
x"3fdc8",
x"3fcad",
x"00353",
x"0031f",
x"3fce1",
x"003ec",
x"3fc14",
x"3fc14",
x"003ec",
x"3fce1",
x"0031f",
x"00353",
x"3fcad",
x"3fdc8",
x"00238",
x"3fc79",
x"00387",
x"003c5",
x"3fc3b",
x"00252",
x"3fdae",
x"3fc2d",
x"003d3",
x"00317",
x"3fce9",
x"00289",
x"3fd77",
x"3fc05",
x"003fb",
x"00322",
x"3fcde",
x"3fcde",
x"00322",
x"003fb",
x"3fc05",
x"3fd77",
x"00289",
x"3fce9",
x"00317",
x"003d3",
x"3fc2d",
x"3fdae",
x"00252",
x"3fc3b",
x"003c5",
x"00387",
x"3fc79",
--Row 28
x"00400",
x"00400",
x"00400",
x"00400",
x"3fc00",
x"3fc00",
x"3fc00",
x"3fc00",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"00000",
x"002d4",
x"002d4",
x"002d4",
x"002d4",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"002d4",
x"002d4",
x"002d4",
x"002d4",
x"3fc4e",
x"3fc4e",
x"3fc4e",
x"3fc4e",
x"003b2",
x"003b2",
x"003b2",
x"003b2",
x"0030f",
x"0030f",
x"0030f",
x"0030f",
x"3fcf1",
x"3fcf1",
x"3fcf1",
x"3fcf1",
x"3fcf1",
x"3fcf1",
x"3fcf1",
x"3fcf1",
x"0030f",
x"0030f",
x"0030f",
x"0030f",
x"003b2",
x"003b2",
x"003b2",
x"003b2",
x"3fc4e",
x"3fc4e",
x"3fc4e",
x"3fc4e",
--Row 29
x"00400",
x"3fc00",
x"00000",
x"00000",
x"3fd2c",
x"002d4",
x"002d4",
x"3fd2c",
x"0030f",
x"3fcf1",
x"003b2",
x"3fc4e",
x"3fc4e",
x"003b2",
x"3fcf1",
x"0030f",
x"00353",
x"3fcad",
x"00238",
x"3fdc8",
x"3fc14",
x"003ec",
x"0031f",
x"3fce1",
x"3fce1",
x"0031f",
x"003ec",
x"3fc14",
x"3fdc8",
x"00238",
x"3fcad",
x"00353",
x"3fc2d",
x"003d3",
x"3fdae",
x"00252",
x"00387",
x"3fc79",
x"3fc3b",
x"003c5",
x"3fcde",
x"00322",
x"3fc05",
x"003fb",
x"00317",
x"3fce9",
x"00289",
x"3fd77",
x"3fd77",
x"00289",
x"3fce9",
x"00317",
x"003fb",
x"3fc05",
x"00322",
x"3fcde",
x"003c5",
x"3fc3b",
x"3fc79",
x"00387",
x"00252",
x"3fdae",
x"003d3",
x"3fc2d",
--Row 30
x"00400",
x"00400",
x"3fc00",
x"3fc00",
x"00000",
x"00000",
x"00000",
x"00000",
x"002d4",
x"002d4",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"3fd2c",
x"002d4",
x"002d4",
x"003b2",
x"003b2",
x"3fc4e",
x"3fc4e",
x"3fcf1",
x"3fcf1",
x"0030f",
x"0030f",
x"0030f",
x"0030f",
x"3fcf1",
x"3fcf1",
x"3fc4e",
x"3fc4e",
x"003b2",
x"003b2",
x"3fc14",
x"3fc14",
x"003ec",
x"003ec",
x"0031f",
x"0031f",
x"3fce1",
x"3fce1",
x"3fdc8",
x"3fdc8",
x"00238",
x"00238",
x"00353",
x"00353",
x"3fcad",
x"3fcad",
x"3fcad",
x"3fcad",
x"00353",
x"00353",
x"00238",
x"00238",
x"3fdc8",
x"3fdc8",
x"3fce1",
x"3fce1",
x"0031f",
x"0031f",
x"003ec",
x"003ec",
x"3fc14",
x"3fc14",
--Row 31
x"00400",
x"3fc00",
x"00000",
x"00000",
x"002d4",
x"3fd2c",
x"3fd2c",
x"002d4",
x"003b2",
x"3fc4e",
x"3fcf1",
x"0030f",
x"0030f",
x"3fcf1",
x"3fc4e",
x"003b2",
x"003ec",
x"3fc14",
x"3fce1",
x"0031f",
x"00238",
x"3fdc8",
x"3fcad",
x"00353",
x"00353",
x"3fcad",
x"3fdc8",
x"00238",
x"0031f",
x"3fce1",
x"3fc14",
x"003ec",
x"3fc05",
x"003fb",
x"00322",
x"3fcde",
x"3fd77",
x"00289",
x"00317",
x"3fce9",
x"3fc79",
x"00387",
x"003c5",
x"3fc3b",
x"3fdae",
x"00252",
x"003d3",
x"3fc2d",
x"3fc2d",
x"003d3",
x"00252",
x"3fdae",
x"3fc3b",
x"003c5",
x"00387",
x"3fc79",
x"3fce9",
x"00317",
x"00289",
x"3fd77",
x"3fcde",
x"00322",
x"003fb",
x"3fc05"
	
);

BEGIN

	indx <= to_integer(unsigned(index));
	coeff <= memory(indx)(WIDTH-1 downto 0);

END dataflow;
